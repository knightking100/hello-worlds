module top;

initial
    $display("Hello, world!");

endmodule
